//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//
// КА с 4мя состояниями. Начальноe состояние при сбросе S0_Idle.
//
// 1) По нажатию кнопки (sync_sw==1 -- сигнал заранее синхронизировали по такту) из начального состояния S0_Idle
// переходим в состояние S1_Wait_1. Если кнопка не нажата, остаёмся в том же состоянии S0_Idle.
// 2) Из состояния S1_Wait_1 переходим в следующее (S2_OK) лишь тогда, когда прождали дребезг(пришёл разрешающий сигнал en==1),
// иначе остаёмся в том же состоянии S1_Wait_1.
// 3) Если находимся в состоянии S2_OK. Если получили сигнал отжатия кнопки (sync_sw==0 -- сигнал заранее синхронизировали по такту),
// то переходим в состояние S3_Wait_2, иначе остаёмся в этом же состоянии S2_OK.
// 4) Из состояния S3_Wait_2 переходим в следующее (S0_Idle) лишь тогда, когда прождали дребезг (пришёл разрешающий сигнал en==1),
// иначе остаёмся в том же состоянии S3_Wait_2.
//
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

module button 
  #(parameter WIDTH_CNT = 24)  // нужно прождать несколько десятков мс в теории, но практика показала, что лучше несколько сотен мс 
  ()                           // подбираем ширину под частоту clk, чтоб отсчитать 100-200 мс
                               // (данная ширина подходит под частоту clk в 100_МГц)

  wire clk;
  reg [WIDTH_CNT-1:0] cnt;  // для хранения пройденного времени от начала нажатия/отжатия кнопки (прожидаем дребезг)
  reg [7:0] cnt_sum;        // количество нажатий кнопки
 

  // состояния State Machine:
  typedef enum reg [1:0]
  { S0_Idle,    // состояние до нажатия кнопки
    S1_Wait_1,  // состояние, когда получен первый импульс нажатой кнопки
    S2_OK,      // состояние, когда прождали дребезг и всё устаканилось
    S3_Wait_2   // состояние, когда получили первый импульс отжатой кнопки
   } st;
 
  st state, next_state;ы
 

  // сигнал, синхронизированный с clk:
  wire sync_sw;
  // синхронизируем нажатие кнопки sw по тактовому сигналу clk и получаем синхронный сигнал sync_sw:
  sync_reg #(1, 0) sync (.clk2(clk), .reset_2(reset_n), .in_clk1(sw), .out_clk2(sync_sw), .kratno(1'b0));
 
 
  always @(posedge clk or negedge reset_n)
    if (!reset_n)
      state <= S0_Idle;
    else
      state <= next_state;

 
  // сигнал ассинхронного сброса счётчика подсчёта времени ожидания
  // (времени, отведённого на дребезг)
  // подсчёт времени ведётся только в состояниях S1_Wait_1 и S3_Wait_2
  wire res_n = !reset_n || ~((state == S1_Wait_1) || (state == S3_Wait_2));  

  // отсчитываем время ожидания до перехода в следующее состояние State Machine (для того, чтоб прождать дребезг)
  always @(posedge clk or posedge res_n)
    if (res_n)
      cnt <= 0;
    else
      cnt <= cnt + 1'b1;
 

  // разрещающий сигнал для перехода в следующее состояние (дребезг прождали)     
  wire en = (cnt[WIDTH_CNT-1]) ? 1 : 0;  // как нужное время прошло, подаём разрешающий сигнал (en=1)

  
  //подсчитываем число нажатий на кнопку: 
  always @(posedge en or negedge reset_n)
    if (!reset_n)
      cnt_sum <= 0;
    else if (state == S1_Wait_1)   // по каждому фронту разрешающего сигнала en, говорящего о том, что дребезг миновал,
      cnt_sum <= cnt_sum + 1'b1;   // и значит, сигнал статичен и соответствует положению кнопки (либо нажата (1), либо отжата (0)) 
                                   // следим за тем, в каком состоянии state мы сейчас находимся.
                            // если мы отсчитали время после нажатия (т.е. state == S1_Wait_1), а не отжатия кнопки, то увеличиваем счётчик числа нажатий
    
  // правила переходов по состояниям: 
  always @*
    case (state)
      S0_Idle   : if (sync_sw)                // Если сейчас S0_Idle, то при условии нажатия на кнопку,
                    next_state = S1_Wait_1;   // переходим в следующее состояние S1_Wait_1;
                  else                        // иначе - 
                    next_state = S0_Idle;     // остаёмся в том же состоянии S0_Idle.
 
      S1_Wait_1 : if (en)                     // Если сейчас S1_Wait_1, то при условии, что уже прождали дребезг,
                    next_state = S2_OK;       // переходим в следующее состояние S2_OK;
                  else                        // иначе -
                    next_state = S1_Wait_1;   // остаёмся в том же состоянии S0_Idle.
 
      S2_OK     : if (!sync_sw)               // Если сейчас S2_OK, то при условии отжатия кнопки,
                    next_state = S3_Wait_2;   // переходим в следующее состояние S3_Wait_2;
                  else                        // иначе - 
                    next_state = S2_OK;       // остаёмся в том же состоянии S2_OK.
                  
      S3_Wait_2 : if (en)                     // Если сейчас S3_Wait_2, то при условии, что уже прождали дребезг,
                    next_state = S0_Idle;     // переходим в следующее состояние S0_Idle;
                  else                        // иначе - 
                    next_state = S3_Wait_2;   // остаёмся в том же состоянии S3_Wait_2.
                             
      default   : next_state = S0_Idle;
 
    endcase
 

  // Если число нажатий на кнопку чётное (в том числе, если не было нажатия), то 1; если нечётное - то 0.
  wire endpoint = (cnt_sum%2) ? 1 : 0; 

endmodule
